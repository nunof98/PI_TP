Circuito com Multiplas Fontes DC (VMalha1 > VMalha2)
V1 1 0 20
V2 3 0 10
R1 1 2 10
R2 2 3 20
R3 2 0 40
.END