Circuito a implementar (Nos impossiveis)
V1 1 3 10
R1 1 3 10
R2 2 0 10
R3 2 0 1
R4 2 3 1
R666 3 1 10
R6 3 0 1
.END