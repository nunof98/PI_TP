Circuito a implementar
V1 1 0 10
R1 1 0 10
R2 2 0 10
R3 2 0 1
R4 2 3 1
R5 2 3 10
R6 3 0 1
.END